-- megafunction wizard: %PLL Reconfig Intel FPGA IP v18.1%
-- GENERATION: XML
-- alt_pll_reconfig.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alt_pll_reconfig is
	generic (
		ENABLE_BYTEENABLE   : boolean := false;
		BYTEENABLE_WIDTH    : integer := 4;
		RECONFIG_ADDR_WIDTH : integer := 6;
		RECONFIG_DATA_WIDTH : integer := 32;
		reconf_width        : integer := 64;
		WAIT_FOR_LOCK       : boolean := true
	);
	port (
		mgmt_clk          : in  std_logic                     := '0';             --          mgmt_clk.clk
		mgmt_reset        : in  std_logic                     := '0';             --        mgmt_reset.reset
		mgmt_waitrequest  : out std_logic;                                        -- mgmt_avalon_slave.waitrequest
		mgmt_read         : in  std_logic                     := '0';             --                  .read
		mgmt_write        : in  std_logic                     := '0';             --                  .write
		mgmt_readdata     : out std_logic_vector(31 downto 0);                    --                  .readdata
		mgmt_address      : in  std_logic_vector(5 downto 0)  := (others => '0'); --                  .address
		mgmt_writedata    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		reconfig_to_pll   : out std_logic_vector(63 downto 0);                    --   reconfig_to_pll.reconfig_to_pll
		reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => '0')  -- reconfig_from_pll.reconfig_from_pll
	);
end entity alt_pll_reconfig;

architecture rtl of alt_pll_reconfig is
	component altera_pll_reconfig_top is
		generic (
			device_family       : string  := "";
			ENABLE_MIF          : boolean := false;
			MIF_FILE_NAME       : string  := "";
			ENABLE_BYTEENABLE   : boolean := false;
			BYTEENABLE_WIDTH    : integer := 4;
			RECONFIG_ADDR_WIDTH : integer := 6;
			RECONFIG_DATA_WIDTH : integer := 32;
			reconf_width        : integer := 64;
			WAIT_FOR_LOCK       : boolean := true
		);
		port (
			mgmt_clk          : in  std_logic                     := 'X';             -- clk
			mgmt_reset        : in  std_logic                     := 'X';             -- reset
			mgmt_waitrequest  : out std_logic;                                        -- waitrequest
			mgmt_read         : in  std_logic                     := 'X';             -- read
			mgmt_write        : in  std_logic                     := 'X';             -- write
			mgmt_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			mgmt_address      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			mgmt_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reconfig_to_pll   : out std_logic_vector(63 downto 0);                    -- reconfig_to_pll
			reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => 'X'); -- reconfig_from_pll
			mgmt_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- byteenable
		);
	end component altera_pll_reconfig_top;

begin

	alt_pll_reconfig_inst : component altera_pll_reconfig_top
		generic map (
			device_family       => "Arria V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => ENABLE_BYTEENABLE,
			BYTEENABLE_WIDTH    => BYTEENABLE_WIDTH,
			RECONFIG_ADDR_WIDTH => RECONFIG_ADDR_WIDTH,
			RECONFIG_DATA_WIDTH => RECONFIG_DATA_WIDTH,
			reconf_width        => reconf_width,
			WAIT_FOR_LOCK       => WAIT_FOR_LOCK
		)
		port map (
			mgmt_clk          => mgmt_clk,          --          mgmt_clk.clk
			mgmt_reset        => mgmt_reset,        --        mgmt_reset.reset
			mgmt_waitrequest  => mgmt_waitrequest,  -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mgmt_read,         --                  .read
			mgmt_write        => mgmt_write,        --                  .write
			mgmt_readdata     => mgmt_readdata,     --                  .readdata
			mgmt_address      => mgmt_address,      --                  .address
			mgmt_writedata    => mgmt_writedata,    --                  .writedata
			reconfig_to_pll   => reconfig_to_pll,   --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => reconfig_from_pll, -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"             --       (terminated)
		);

end architecture rtl; -- of alt_pll_reconfig
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2024 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_pll_reconfig" version="18.1" >
-- Retrieval info: 	<generic name="device_family" value="Arria V" />
-- Retrieval info: 	<generic name="ENABLE_MIF" value="false" />
-- Retrieval info: 	<generic name="MIF_FILE_NAME" value="" />
-- Retrieval info: 	<generic name="ENABLE_BYTEENABLE" value="false" />
-- Retrieval info: </instance>
-- IPFS_FILES : alt_pll_reconfig.vho
-- RELATED_FILES: alt_pll_reconfig.vhd, altera_pll_reconfig_top.v, altera_pll_reconfig_core.v, altera_std_synchronizer.v
